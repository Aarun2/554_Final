module fetch_buffer();
  
  
endmodule

module br_predict();
  
  
endmodule

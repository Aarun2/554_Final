module buffer();
  input [size-1:0] instr;
  
endmodule
